*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Wed Oct 24 2018 at 13:40:17

*
* Globals.
*
.global VSS VDD


*
* Component pathname : $MGC_DESIGN_KIT/symbols/ncap [SPICE]
*
*       .include /mgc/v9.0d_rhelx86linux/icstation_home/mgc_icstd_lib/mit0.25/symbols/ncap/NCAP

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/HW6/npcmos_hw6
*
        X1 F VSS VSS NCAP CAPACITANCE=20F
        V1 VDD VSS DC 2.5V
        M8 F CLK_NOT VSS VSS NMOS L=1.2u W=2.4u M=1
        M7 F C_NOT N$12 VDD PMOS L=2.0u W=400.0u M=1
        M6 F A N$37 VDD PMOS L=2.0u W=20.0u M=1
        M5 N$37 N$10 N$12 VDD PMOS L=2.0u W=20.0u M=1
        M4 N$35 CLK VSS VSS NMOS L=1.2u W=2.4u M=1
        M3 N$12 CLK_NOT VDD VDD PMOS L=2.0u W=30.0u M=1
        M2 N$10 B N$35 VSS NMOS L=1.2u W=2.4u M=1
        M1 N$10 CLK VDD VDD PMOS L=2.0u W=30.0u M=1
*
.end
