* Component: /home/ece_lab/mentor/ECE4500/Lab7/two_input_nand  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/Lab7/two_input_nand/eldonet/two_input_nand_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 400N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A_NOT) V(B) V(B_NOT) V(F)

* --- Params
.TEMP 27

* --- Forces
VFORCE__T A_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0011 R
VFORCE__T_1 B VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0101 R
VFORCE__T_2 B_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1010 R

* --- Libsetup

