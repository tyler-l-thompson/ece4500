* Component: /home/ece_lab/mentor/ECE4500/Project1/full_add_sub  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/Project1/full_add_sub/eldonet/full_add_sub_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 3200N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A) V(A_NOT) V(A_XOR_B) V(A_XOR_B_NOT) V(BIN_CIN) V(BOUT_COUT)
+ V(CC0) V(CC0_NOT) V(CC3) V(CC3_NOT)
.PROBE TRAN V(SUM_D)

* --- Params
.TEMP 27

* --- Forces
VFORCE__Bin_Cin BIN_CIN VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 01010101010101010101010101010101 R
VFORCE__CC0 CC0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 00000000111111110000000011111111 R
VFORCE__CC0_not CC0_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 11111111000000001111111100000000 R
VFORCE__CC3 CC3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 000000000000000011111111111111111 R
VFORCE__CC3_not CC3_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 111111111111111110000000000000000 R
VFORCE__A_xor_B A_XOR_B VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 00111100001111000011110000111100 R
VFORCE__A_xor_B_not A_XOR_B_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 11000011110000111100001111000011 R
VFORCE__A_not_1 A_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 11110000111100001111000011110000 R
VFORCE__A A VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 00001111000011110000111100001111 R

* --- Libsetup

