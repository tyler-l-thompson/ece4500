*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Fri Oct 19 2018 at 02:28:38

*
* Globals.
*
.global VSS VDD

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/Project1/two_input_mux/two_input_mux
*
        V1 VDD VSS DC 2.5V
        M4 F SELECT A VSS NMOS L=1.2u W=2.4u M=1
        M3 F SELECT_NOT A VDD PMOS L=1.2u W=2.4u M=1
        M2 F SELECT_NOT B VSS NMOS L=1.2u W=2.4u M=1
        M1 F SELECT B VDD PMOS L=1.2u W=2.4u M=1
*
.end
