*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Sat Oct 27 2018 at 11:22:27

*
* Globals.
*
.global VDD VSS

*
* Component pathname : /home/ece_lab/mentor/4500/Project_1/4input_MUX
*
.subckt 4INPUT_MUX  F0 F1 F2 F3 A0 A1 A2 A3 B0 B1 B2 B3 SEL SEL_NOT

        M16 B3 SEL F3 VSS NMOS L=1.2u W=2u M=1
        M15 B3 SEL_NOT F3 VDD PMOS L=1.2u W=7.5u M=1
        M14 A3 SEL_NOT F3 VSS NMOS L=1.2u W=2u M=1
        M13 A3 SEL F3 VDD PMOS L=1.2u W=7.5u M=1
        M12 B2 SEL F2 VSS NMOS L=1.2u W=2u M=1
        M11 B2 SEL_NOT F2 VDD PMOS L=1.2u W=7.5u M=1
        M10 A2 SEL_NOT F2 VSS NMOS L=1.2u W=2u M=1
        M9 A2 SEL F2 VDD PMOS L=1.2u W=7.5u M=1
        M8 B1 SEL F1 VSS NMOS L=1.2u W=2u M=1
        M7 B1 SEL_NOT F1 VDD PMOS L=1.2u W=7.5u M=1
        M6 A1 SEL_NOT F1 VSS NMOS L=1.2u W=2u M=1
        M5 A1 SEL F1 VDD PMOS L=1.2u W=7.5u M=1
        M4 B0 SEL F0 VSS NMOS L=1.2u W=2u M=1
        M3 B0 SEL_NOT F0 VDD PMOS L=1.2u W=7.5u M=1
        M2 A0 SEL_NOT F0 VSS NMOS L=1.2u W=2u M=1
        M1 A0 SEL F0 VDD PMOS L=1.2u W=7.5u M=1
.ends 4INPUT_MUX

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/4500/Project_1/Project_1_MUX
*
        X_4INPUT_MUX7 N$53 N$55 N$57 N$59 ZERO0 ZERO1 ZERO2 ZERO3 A_PLUS_B_WITH_CARRY0
+ A_PLUS_B_WITH_CARRY1 A_PLUS_B_WITH_CARRY2 A_PLUS_B_WITH_CARRY3 CC0 CC0_NOT 4INPUT_MUX
        X_4INPUT_MUX6 N$45 N$47 N$49 N$51 ASLA0 ASLA1 ASLA2 ASLA3 ASRA0
+ ASRA1 ASRA2 ASRA3 CC0 CC0_NOT 4INPUT_MUX
        V1 VDD VSS DC 2.5V
        X_4INPUT_MUX15 F0 F1 F2 F3 N$101 N$103 N$105 N$109 N$288 N$289 N$290
+ N$291 CC3 CC3_NOT 4INPUT_MUX
        X_4INPUT_MUX14 N$288 N$289 N$290 N$291 N$69 N$71 N$73 N$75 N$77
+ N$79 N$81 N$83 CC2 CC2_NOT 4INPUT_MUX
        X_4INPUT_MUX13 N$101 N$103 N$105 N$109 N$85 N$87 N$89 N$91 N$93
+ N$95 N$97 N$99 CC2 CC2_NOT 4INPUT_MUX
        X_4INPUT_MUX12 N$77 N$79 N$81 N$83 N$53 N$55 N$57 N$59 N$61 N$63
+ N$65 N$67 CC1 CC1_NOT 4INPUT_MUX
        X_4INPUT_MUX11 N$69 N$71 N$73 N$75 N$36 N$38 N$39 N$41 N$45 N$47
+ N$49 N$51 CC1 CC1_NOT 4INPUT_MUX
        X_4INPUT_MUX10 N$93 N$95 N$97 N$99 N$20 N$22 N$24 N$25 N$27 N$29
+ N$31 N$33 CC1 CC1_NOT 4INPUT_MUX
        X_4INPUT_MUX9 N$85 N$87 N$89 N$91 N$2 N$4 N$9 N$8 N$12 N$14 N$16
+ N$18 CC1 CC1_NOT 4INPUT_MUX
        X_4INPUT_MUX8 N$61 N$63 N$65 N$67 A_MINUS_B_WITH_BORROW0 A_MINUS_B_WITH_BORROW1
+ A_MINUS_B_WITH_BORROW2 A_MINUS_B_WITH_BORROW3 B_PLUS_ONE0 B_PLUS_ONE1
+ B_PLUS_ONE2 B_PLUS_ONE3 CC0 CC0_NOT 4INPUT_MUX
        X_4INPUT_MUX5 N$36 N$38 N$39 N$41 LSLA0 LSLA1 LSLA2 LSLA3 LSRA0
+ LSRA1 LSRA2 LSRA3 CC0 CC0_NOT 4INPUT_MUX
        X_4INPUT_MUX4 N$27 N$29 N$31 N$33 A_MINUS_B0 A_MINUS_B1 A_MINUS_B2
+ A_MINUS_B3 B0 B1 B2 B3 CC0 CC0_NOT 4INPUT_MUX
        X_4INPUT_MUX3 N$20 N$22 N$24 N$25 A_XOR_B0 A_XOR_B1 A_XOR_B2 A_XOR_B3
+ A_PLUS_B0 A_PLUS_B1 A_PLUS_B2 A_PLUS_B3 CC0 CC0_NOT 4INPUT_MUX
        X_4INPUT_MUX2 N$12 N$14 N$16 N$18 A_AND_B0 A_AND_B1 A_AND_B2 A_AND_B3
+ A_OR_B0 A_OR_B1 A_OR_B2 A_OR_B3 CC0 CC0_NOT 4INPUT_MUX
        X_4INPUT_MUX1 N$2 N$4 N$9 N$8 A0 A1 A2 A3 A0_NOT A1_NOT A2_NOT A3_NOT
+ CC0 CC0_NOT 4INPUT_MUX
*
.end
