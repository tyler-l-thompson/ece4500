*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Tue Oct 30 2018 at 11:53:38

*
* Globals.
*
.global VDD VSS

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/one_input_inverter/one_input_inverter
*
.subckt ONE_INPUT_INVERTER  OUT IN VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        M2 OUT IN VSS VSS NMOS L=1.2u W=2.25u M=1
        M1 OUT IN VDD VDD PMOS L=1.2u W=6.75u M=1
.ends ONE_INPUT_INVERTER

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/Lab8/3_state_buffer/3_state_buffer
*
        V1 VDD VSS DC 2.5V
        X_ONE_INPUT_INVERTER1 N$17 DOUT_18 VDD VSS ONE_INPUT_INVERTER
        M4 N$19 N$17 VDD VDD PMOS L=1.2u W=13.5u M=1
        M3 DOUTB_18 DEN_NOT_18 N$19 VDD PMOS L=1.2u W=13.5u M=1
        M2 DOUTB_18 DEN_18 N$4 VSS NMOS L=1.2u W=4.8u M=1
        M1 N$4 N$17 VSS VSS NMOS L=1.2u W=4.8u M=1
*
.end
