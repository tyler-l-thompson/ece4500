*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Tue Oct 23 2018 at 20:34:45

*
* Globals.
*
.global VDD VSS

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/one_input_inverter/one_input_inverter
*
.subckt ONE_INPUT_INVERTER  OUT IN VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        M2 OUT IN VSS VSS NMOS L=1.2u W=2.25u M=1
        M1 OUT IN VDD VDD PMOS L=1.2u W=6.75u M=1
.ends ONE_INPUT_INVERTER

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Lab7/two_input_and
*
.subckt TWO_INPUT_AND  F A B VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        M4 A N$15 F VDD PMOS L=1.2u W=2.4u M=1
        M3 A B F VSS NMOS L=1.2u W=2.4u M=1
        X_ONE_INPUT_INVERTER1 N$15 B VDD VSS ONE_INPUT_INVERTER
        M2 F N$15 B VSS NMOS L=1.2u W=2.4u M=1
        M1 A B F VSS NMOS L=1.2u W=2.4u M=1
.ends TWO_INPUT_AND

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Lab7/three_input_and
*
.subckt THREE_INPUT_AND  F A B C VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        X_TWO_INPUT_AND2 F N$46 C VDD VSS TWO_INPUT_AND
        X_TWO_INPUT_AND1 N$46 A B VDD VSS TWO_INPUT_AND
.ends THREE_INPUT_AND

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Lab7/asynchronous_sr_latch
*
.subckt ASYNCHRONOUS_SR_LATCH  QN_18 QN_NOT_18 CLR_NOT_18 R_18 S_18 VDD_ESC1
+ VSS_ESC2

        .CONNECT VDD VDD_ESC1
        .CONNECT VSS VSS_ESC2
        M7 QN_18 R_18 VSS VSS NMOS L=2.0u W=12.0u M=1
        M1 QN_18 CLR_NOT_18 VSS VSS NMOS L=2.0u W=12.0u M=1
        M8 QN_NOT_18 S_18 VSS VSS NMOS L=2.0u W=12.0u M=1
        M5 QN_NOT_18 QN_18 VSS VSS NMOS L=2.0u W=3.0u M=1
        M4 QN_18 QN_NOT_18 VSS VSS NMOS L=2.0u W=3.0u M=1
        M3 QN_NOT_18 QN_18 VDD VDD PMOS L=2.0u W=9.0u M=1
        M2 QN_18 QN_NOT_18 VDD VDD PMOS L=2.0u W=9.0u M=1
.ends ASYNCHRONOUS_SR_LATCH

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Lab7/two_input_nor
*
.subckt TWO_INPUT_NOR  F A_NOT B B_NOT VDD_ESC1

        .CONNECT VDD VDD_ESC1
        M5 A_NOT B F VDD PMOS L=1.2u W=2.4u M=1
        M3 A_NOT B_NOT F VSS NMOS L=1.2u W=2.4u M=1
        M2 F B B_NOT VSS NMOS L=1.2u W=2.4u M=1
        M1 A_NOT B_NOT F VSS NMOS L=1.2u W=2.4u M=1
.ends TWO_INPUT_NOR

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Lab7/t_flip_flop
*
.subckt T_FLIP_FLOP  QN_18 QN_NOT_18 CLK_18 CLR_NOT_18 T_18 VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        X_ONE_INPUT_INVERTER24 N$432 N$407 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER23 N$407 N$416 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER22 N$431 N$401 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER21 N$401 N$415 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER2 N$313 N$427 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER1 N$357 N$296 VDD VSS ONE_INPUT_INVERTER
        X_THREE_INPUT_AND2 N$302 CLK_18 T_18 QN_NOT_18 VDD VSS THREE_INPUT_AND
        X_THREE_INPUT_AND1 N$296 CLK_18 T_18 QN_18 VDD VSS THREE_INPUT_AND
        X_ONE_INPUT_INVERTER3 N$189 CLR_NOT_18 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER18 N$415 N$385 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER17 N$385 N$399 VDD VSS ONE_INPUT_INVERTER
        X_ASYNCHRONOUS_SR_LATCH1 QN_18 QN_NOT_18 N$189 N$337 N$336 VDD VSS ASYNCHRONOUS_SR_LATCH
        X_ONE_INPUT_INVERTER14 N$399 N$364 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER13 N$364 N$378 VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_NOR2 N$336 N$330 N$334 N$321 VDD TWO_INPUT_NOR
        X_TWO_INPUT_NOR1 N$337 N$330 N$314 N$313 VDD TWO_INPUT_NOR
        X_ONE_INPUT_INVERTER7 N$334 N$321 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER4 N$314 N$313 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER9 N$354 N$351 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER10 N$378 N$354 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER26 N$421 N$418 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER25 N$418 N$431 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER8 N$330 CLK_18 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER16 N$400 N$370 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER15 N$370 N$379 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER12 N$379 N$360 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER11 N$360 N$357 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER6 N$321 N$421 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER5 N$351 N$302 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER20 N$416 N$391 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER19 N$391 N$400 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER28 N$427 N$424 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER27 N$424 N$432 VDD VSS ONE_INPUT_INVERTER
.ends T_FLIP_FLOP

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/Lab7/three_bit_synchronous_counter
*
        X_TWO_INPUT_AND4 CY_18 N$147 N$150 VDD VSS TWO_INPUT_AND
        X_TWO_INPUT_AND3 N$150 Q2_18 CLK_18 VDD VSS TWO_INPUT_AND
        X_TWO_INPUT_AND2 N$147 Q0_18 Q1_18 VDD VSS TWO_INPUT_AND
        X_TWO_INPUT_AND1 N$143 Q0_18 Q1_18 VDD VSS TWO_INPUT_AND
        X_T_FLIP_FLOP3 Q2_18 N$89 CLK_18 CLR_NOT_18 N$143 VDD VSS T_FLIP_FLOP
        X_T_FLIP_FLOP2 Q1_18 N$87 CLK_18 CLR_NOT_18 Q0_18 VDD VSS T_FLIP_FLOP
        X_T_FLIP_FLOP1 Q0_18 N$84 CLK_18 CLR_NOT_18 VDD VDD VSS T_FLIP_FLOP
        V1 VDD VSS DC 2.5V
*
.end
