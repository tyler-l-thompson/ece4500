*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Fri Oct 19 2018 at 16:47:44

*
* Globals.
*
.global VSS VDD

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/Project1/two_input_and/two_input_and
*
        V1 VDD VSS DC 2.5V
        M4 F B_NOT VSS VSS NMOS L=1.2u W=2.4u M=1
        M3 F A_NOT VSS VSS NMOS L=1.2u W=2.4u M=1
        M2 F B_NOT N$17 VDD PMOS L=1.2u W=2.4u M=1
        M1 N$17 A_NOT VDD VDD PMOS L=1.2u W=2.4u M=1
*
.end
