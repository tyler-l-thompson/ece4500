*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Sun Oct 28 2018 at 06:46:53

*
* Globals.
*
.global VDD VSS

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/one_input_inverter/one_input_inverter
*
.subckt ONE_INPUT_INVERTER  OUT IN VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        M2 OUT IN VSS VSS NMOS L=1.2u W=2.25u M=1
        M1 OUT IN VDD VDD PMOS L=1.2u W=6.75u M=1
.ends ONE_INPUT_INVERTER

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/two_input_and_2/two_input_and
*
.subckt TWO_INPUT_AND  F A B B_NOT VDD_ESC1

        .CONNECT VDD VDD_ESC1
        M5 A B F VSS NMOS L=1.2u W=2.4u M=1
        M4 F B_NOT B VSS NMOS L=1.2u W=2.4u M=1
        M3 A B F VSS NMOS L=1.2u W=2.4u M=1
        M2 A B_NOT F VDD PMOS L=1.2u W=2.4u M=1
.ends TWO_INPUT_AND

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/add_sub_ovf_sel/add_sub_ovf_sel
*
.subckt ADD_SUB_OVF_SEL  F CC0 CC0_NOT CC1 CC1_NOT CC2_NOT CC3_NOT VDD_ESC1
+ VSS_ESC2

        .CONNECT VDD VDD_ESC1
        .CONNECT VSS VSS_ESC2
        M8 N$28 CC0 N$24 VDD PMOS L=1.2u W=5.0u M=1
        M18 N$50 CC1_NOT VSS VSS NMOS L=1.2u W=2.4u M=1
        M17 N$50 CC2_NOT VSS VSS NMOS L=1.2u W=2.4u M=1
        M16 N$50 CC0 VSS VSS NMOS L=1.2u W=2.4u M=1
        M15 N$41 CC3_NOT N$50 VSS NMOS L=1.2u W=2.4u M=1
        M14 N$41 CC2_NOT N$50 VSS NMOS L=1.2u W=2.4u M=1
        M13 N$41 CC0_NOT N$50 VSS NMOS L=1.2u W=2.4u M=1
        M12 F CC1 N$41 VSS NMOS L=1.2u W=2.4u M=1
        M11 F CC2_NOT N$41 VSS NMOS L=1.2u W=2.4u M=1
        M10 F CC0_NOT N$41 VSS NMOS L=1.2u W=2.4u M=1
        M9 F CC1_NOT N$28 VDD PMOS L=1.2u W=5.0u M=1
        M7 N$24 CC2_NOT VDD VDD PMOS L=1.2u W=5.0u M=1
        M6 F CC0_NOT N$18 VDD PMOS L=1.2u W=5.0u M=1
        M5 N$18 CC3_NOT N$14 VDD PMOS L=1.2u W=5.0u M=1
        M4 N$14 CC2_NOT VDD VDD PMOS L=1.2u W=5.0u M=1
        M3 F CC2_NOT N$12 VDD PMOS L=1.2u W=5.0u M=1
        M2 N$12 CC1 N$8 VDD PMOS L=1.2u W=5.0u M=1
        M1 N$8 CC0_NOT VDD VDD PMOS L=1.2u W=5.0u M=1
.ends ADD_SUB_OVF_SEL

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/one_input_buffer/one_input_buffer
*
.subckt ONE_INPUT_BUFFER  OUT IN VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        X_ONE_INPUT_INVERTER2 OUT N$3 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER1 N$3 IN VDD VSS ONE_INPUT_INVERTER
.ends ONE_INPUT_BUFFER

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/two_input_xor/two_input_xor
*
.subckt TWO_INPUT_XOR  F A A_NOT B VDD_ESC1

        .CONNECT VDD VDD_ESC1
        M4 F A_NOT B VSS NMOS L=1.2u W=2.4u M=1
        M3 F A B VDD PMOS L=1.2u W=2.4u M=1
        M2 F B A_NOT VSS NMOS L=1.2u W=2.4u M=1
        M1 F B A VDD PMOS L=1.2u W=2.4u M=1
.ends TWO_INPUT_XOR

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/two_input_mux/two_input_mux
*
.subckt TWO_INPUT_MUX  F A B SELECT SELECT_NOT VDD_ESC1

        .CONNECT VDD VDD_ESC1
        M4 F SELECT B VDD PMOS L=1.2u W=2.4u M=1
        M3 F SELECT_NOT B VSS NMOS L=1.2u W=2.4u M=1
        M2 F SELECT_NOT A VDD PMOS L=1.2u W=2.4u M=1
        M1 F SELECT A VSS NMOS L=1.2u W=2.4u M=1
.ends TWO_INPUT_MUX

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/two_input_or/two_input_or
*
.subckt TWO_INPUT_OR  F A_NOT B_NOT VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        M3 N$11 B_NOT VSS VSS NMOS L=1.2u W=6.4u M=1
        M2 F A_NOT N$11 VSS NMOS L=1.2u W=6.4u M=1
        M1 F VSS VDD VDD PMOS L=4.8u W=2.4u M=1
.ends TWO_INPUT_OR

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/full_add_sub/full_add_sub
*
.subckt FULL_ADD_SUB  BOUT_COUT SUM_DIFF A A_NOT A_XOR_B A_XOR_B_NOT BIN_CIN
+ CC0 CC0_NOT CC3 CC3_NOT VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        X_TWO_INPUT_XOR1 SUM_DIFF A_XOR_B A_XOR_B_NOT N$39 VDD TWO_INPUT_XOR
        X_TWO_INPUT_MUX4 N$39 BIN_CIN VSS CC3 CC3_NOT VDD TWO_INPUT_MUX
        X_TWO_INPUT_MUX3 BOUT_COUT N$11 N$9 CC0 CC0_NOT VDD TWO_INPUT_MUX
        X_TWO_INPUT_MUX2 N$9 A_NOT N$39 A_XOR_B A_XOR_B_NOT VDD TWO_INPUT_MUX
        X_TWO_INPUT_MUX1 N$11 N$39 A A_XOR_B A_XOR_B_NOT VDD TWO_INPUT_MUX
.ends FULL_ADD_SUB

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/one_bit_alu/one_bit_alu
*
.subckt ONE_BIT_ALU  A_AND_B A_NOT A_OR_B A_XOR_B BOUT_COUT SUM_DIFF A ADD
+ B BIN_CIN CC0 CC0_NOT CC1 CC1_NOT CC3 CC3_NOT VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        X_TWO_INPUT_MUX2 N$129 N$130 A CC0 CC0_NOT VDD TWO_INPUT_MUX
        X_TWO_INPUT_OR1 A_OR_B A_NOT N$10 VDD VSS TWO_INPUT_OR
        X_TWO_INPUT_MUX1 N$130 ADD A N$142 N$143 VDD TWO_INPUT_MUX
        X_ONE_INPUT_INVERTER3 N$10 B VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER2 A_NOT A VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_AND1 A_AND_B A B N$10 VDD TWO_INPUT_AND
        X_ONE_INPUT_INVERTER1 N$22 A_XOR_B VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_XOR1 A_XOR_B B N$10 N$129 VDD TWO_INPUT_XOR
        X_ONE_INPUT_INVERTER5 N$143 N$142 VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_AND2 N$142 CC0 CC1 CC1_NOT VDD TWO_INPUT_AND
        X_FULL_ADD_SUB1 BOUT_COUT SUM_DIFF N$130 N$122 A_XOR_B N$22 BIN_CIN
+ CC0 CC0_NOT CC3 CC3_NOT VDD VSS FULL_ADD_SUB
        X_ONE_INPUT_INVERTER4 N$122 N$129 VDD VSS ONE_INPUT_INVERTER
.ends ONE_BIT_ALU

*
* Component pathname : /home/ece_lab/mentor/ECE4500/Project1/four_input_and/four_input_and
*
.subckt FOUR_INPUT_AND  F A B B_NOT C D D_NOT VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        X_ONE_INPUT_INVERTER1 N$4 N$5 VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_AND3 F N$7 N$5 N$4 VDD TWO_INPUT_AND
        X_TWO_INPUT_AND2 N$5 C D D_NOT VDD TWO_INPUT_AND
        X_TWO_INPUT_AND1 N$7 A B B_NOT VDD TWO_INPUT_AND
.ends FOUR_INPUT_AND

*
* Component pathname : /home/ece_lab/mentor/4500/Project_1/4input_MUX
*
.subckt 4INPUT_MUX  F0 F1 F2 F3 A0 A1 A2 A3 B0 B1 B2 B3 SEL SEL_NOT VDD_ESC1

        .CONNECT VDD VDD_ESC1
        M16 B3 SEL F3 VSS NMOS L=1.2u W=2u M=1
        M15 B3 SEL_NOT F3 VDD PMOS L=1.2u W=7.5u M=1
        M14 A3 SEL_NOT F3 VSS NMOS L=1.2u W=2u M=1
        M13 A3 SEL F3 VDD PMOS L=1.2u W=7.5u M=1
        M12 B2 SEL F2 VSS NMOS L=1.2u W=2u M=1
        M11 B2 SEL_NOT F2 VDD PMOS L=1.2u W=7.5u M=1
        M10 A2 SEL_NOT F2 VSS NMOS L=1.2u W=2u M=1
        M9 A2 SEL F2 VDD PMOS L=1.2u W=7.5u M=1
        M8 B1 SEL F1 VSS NMOS L=1.2u W=2u M=1
        M7 B1 SEL_NOT F1 VDD PMOS L=1.2u W=7.5u M=1
        M6 A1 SEL_NOT F1 VSS NMOS L=1.2u W=2u M=1
        M5 A1 SEL F1 VDD PMOS L=1.2u W=7.5u M=1
        M4 B0 SEL F0 VSS NMOS L=1.2u W=2u M=1
        M3 B0 SEL_NOT F0 VDD PMOS L=1.2u W=7.5u M=1
        M2 A0 SEL_NOT F0 VSS NMOS L=1.2u W=2u M=1
        M1 A0 SEL F0 VDD PMOS L=1.2u W=7.5u M=1
.ends 4INPUT_MUX

*
* Component pathname : /home/ece_lab/mentor/4500/Project_1/Project_1_MUX
*
.subckt PROJECT_1_MUX  F0 F1 F2 F3 A0 A0_NOT A1 A1_NOT A2 A2_NOT A3 A3_NOT
+ A_AND_B0 A_AND_B1 A_AND_B2 A_AND_B3 A_MINUS_B0 A_MINUS_B1 A_MINUS_B2 A_MINUS_B3
+ A_MINUS_B_WITH_BORROW0 A_MINUS_B_WITH_BORROW1 A_MINUS_B_WITH_BORROW2 A_MINUS_B_WITH_BORROW3
+ A_OR_B0 A_OR_B1 A_OR_B2 A_OR_B3 A_PLUS_B0 A_PLUS_B1 A_PLUS_B2 A_PLUS_B3
+ A_PLUS_B_WITH_CARRY0 A_PLUS_B_WITH_CARRY1 A_PLUS_B_WITH_CARRY2 A_PLUS_B_WITH_CARRY3
+ A_XOR_B0 A_XOR_B1 A_XOR_B2 A_XOR_B3 ASLA0 ASLA1 ASLA2 ASLA3 ASRA0 ASRA1
+ ASRA2 ASRA3 B0 B1 B2 B3 B_PLUS_ONE0 B_PLUS_ONE1 B_PLUS_ONE2 B_PLUS_ONE3
+ CC0 CC0_NOT CC1 CC1_NOT CC2 CC2_NOT CC3 CC3_NOT LSLA0 LSLA1 LSLA2 LSLA3
+ LSRA0 LSRA1 LSRA2 LSRA3 VDD_ESC1 ZERO0 ZERO1 ZERO2 ZERO3

        .CONNECT VDD VDD_ESC1
        X_4INPUT_MUX6 N$45 N$47 N$49 N$51 ASLA0 ASLA1 ASLA2 ASLA3 ASRA0
+ ASRA1 ASRA2 ASRA3 CC0 CC0_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX5 N$36 N$38 N$39 N$41 LSLA0 LSLA1 LSLA2 LSLA3 LSRA0
+ LSRA1 LSRA2 LSRA3 CC0 CC0_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX4 N$27 N$29 N$31 N$33 A_MINUS_B0 A_MINUS_B1 A_MINUS_B2
+ A_MINUS_B3 B0 B1 B2 B3 CC0 CC0_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX3 N$20 N$22 N$24 N$25 A_XOR_B0 A_XOR_B1 A_XOR_B2 A_XOR_B3
+ A_PLUS_B0 A_PLUS_B1 A_PLUS_B2 A_PLUS_B3 CC0 CC0_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX2 N$12 N$14 N$16 N$18 A_AND_B0 A_AND_B1 A_AND_B2 A_AND_B3
+ A_OR_B0 A_OR_B1 A_OR_B2 A_OR_B3 CC0 CC0_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX1 N$2 N$4 N$9 N$8 A0 A1 A2 A3 A0_NOT A1_NOT A2_NOT A3_NOT
+ CC0 CC0_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX13 N$101 N$103 N$105 N$109 N$85 N$87 N$89 N$91 N$93
+ N$95 N$97 N$99 CC2 CC2_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX12 N$85 N$87 N$89 N$91 N$2 N$4 N$9 N$8 N$12 N$14 N$16
+ N$18 CC1 CC1_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX11 N$93 N$95 N$97 N$99 N$20 N$22 N$24 N$25 N$27 N$29
+ N$31 N$33 CC1 CC1_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX10 N$69 N$71 N$73 N$75 N$36 N$38 N$39 N$41 N$45 N$47
+ N$49 N$51 CC1 CC1_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX9 N$77 N$79 N$81 N$83 N$53 N$55 N$57 N$59 N$61 N$63
+ N$65 N$67 CC1 CC1_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX8 N$61 N$63 N$65 N$67 A_MINUS_B_WITH_BORROW0 A_MINUS_B_WITH_BORROW1
+ A_MINUS_B_WITH_BORROW2 A_MINUS_B_WITH_BORROW3 B_PLUS_ONE0 B_PLUS_ONE1
+ B_PLUS_ONE2 B_PLUS_ONE3 CC0 CC0_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX7 N$53 N$55 N$57 N$59 ZERO0 ZERO1 ZERO2 ZERO3 A_PLUS_B_WITH_CARRY0
+ A_PLUS_B_WITH_CARRY1 A_PLUS_B_WITH_CARRY2 A_PLUS_B_WITH_CARRY3 CC0 CC0_NOT
+ VDD 4INPUT_MUX
        X_4INPUT_MUX14 N$288 N$289 N$290 N$291 N$69 N$71 N$73 N$75 N$77
+ N$79 N$81 N$83 CC2 CC2_NOT VDD 4INPUT_MUX
        X_4INPUT_MUX15 F0 F1 F2 F3 N$101 N$103 N$105 N$109 N$288 N$289 N$290
+ N$291 CC3 CC3_NOT VDD 4INPUT_MUX
.ends PROJECT_1_MUX

*
* Component pathname : /home/ece_lab/mentor/4500/Project_1/Shifts
*
.subckt SHIFTS  F0 F1 F2 F3 OVF A0 A1 A2 A3 C_OUT CC0 CC0_NOT CC1 CC1_NOT
+ VDD_ESC1 VSS_ESC2

        .CONNECT VSS VSS_ESC2
        .CONNECT VDD VDD_ESC1
        M5 A2 CC0 F3 VDD PMOS L=1.2u W=7.5u M=1
        M3 A3 CC1_NOT C_OUT VDD PMOS L=1.2u W=7.5u M=1
        M4 A3 CC1 C_OUT VSS NMOS L=1.2u W=2u M=1
        M1 VSS CC1 C_OUT VDD PMOS L=1.2u W=7.5u M=1
        M2 VSS CC1_NOT C_OUT VSS NMOS L=1.2u W=2u M=1
        M20 A1 CC0 F0 VSS NMOS L=1.2u W=2u M=1
        M18 VSS CC0_NOT F0 VSS NMOS L=1.2u W=2u M=1
        M19 A1 CC0_NOT F0 VDD PMOS L=1.2u W=7.5u M=1
        M21 C_OUT CC0 OVF VDD PMOS L=1.2u W=7.5u M=1
        M24 VSS CC0 OVF VSS NMOS L=1.2u W=2u M=1
        M23 VSS CC0_NOT OVF VDD PMOS L=1.2u W=7.5u M=1
        M22 C_OUT CC0_NOT OVF VSS NMOS L=1.2u W=2u M=1
        M6 A2 CC0_NOT F3 VSS NMOS L=1.2u W=2u M=1
        M17 VSS CC0 F0 VDD PMOS L=1.2u W=7.5u M=1
        M16 A2 CC0 F1 VSS NMOS L=1.2u W=2u M=1
        M15 A2 CC0_NOT F1 VDD PMOS L=1.2u W=7.5u M=1
        M14 A0 CC0_NOT F1 VSS NMOS L=1.2u W=2u M=1
        M13 A0 CC0 F1 VDD PMOS L=1.2u W=7.5u M=1
        M12 A3 CC0 F2 VSS NMOS L=1.2u W=2u M=1
        M11 A3 CC0_NOT F2 VDD PMOS L=1.2u W=7.5u M=1
        M10 A1 CC0_NOT F2 VSS NMOS L=1.2u W=2u M=1
        M9 A1 CC0 F2 VDD PMOS L=1.2u W=7.5u M=1
        M8 C_OUT CC0 F3 VSS NMOS L=1.2u W=2u M=1
        M7 C_OUT CC0_NOT F3 VDD PMOS L=1.2u W=7.5u M=1
.ends SHIFTS

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/Project1/four_bit_alu/four_bit_alu
*
        V1 VDD VSS DC 2.5V
        X_ONE_INPUT_INVERTER11 N$492 OVF_SEL1 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER5 N$115 N$103 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER6 N$119 N$118 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER7 N$123 N$282 VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_AND1 OVF_SEL1 CC3 N$555 CC2 VDD TWO_INPUT_AND
        X_ONE_INPUT_INVERTER2 N$555 CC2 VDD VSS ONE_INPUT_INVERTER
        X_ADD_SUB_OVF_SEL1 OVF_SEL0 CC0 N$583 CC1 N$629 N$555 N$553 VDD
+ VSS ADD_SUB_OVF_SEL
        X_ONE_INPUT_BUFFER9 OVF N$475 VDD VSS ONE_INPUT_BUFFER
        X_ONE_INPUT_BUFFER8 Z N$615 VDD VSS ONE_INPUT_BUFFER
        X_TWO_INPUT_XOR1 ADD_OVF N$369 N$367 COUT_2 VDD TWO_INPUT_XOR
        X_I$3 N$30 N$31 N$32 N$33 COUT_1 N$36 A1 VSS B1 COUT_0 CC0 N$583
+ CC1 N$629 VDD VSS VDD VSS ONE_BIT_ALU
        X_I$2 N$19 N$20 N$21 A_XOR_B_2 N$369 N$26 A3 VSS B3 COUT_2 CC0 N$583
+ CC1 N$629 VDD VSS VDD VSS ONE_BIT_ALU
        X_I$1 N$65 N$66 N$67 N$68 N$568 N$70 A2 VSS B2 COUT_1 CC0 N$583
+ CC1 N$629 VDD VSS VDD VSS ONE_BIT_ALU
        X_ONE_INPUT_BUFFER1 S N$282 VDD VSS ONE_INPUT_BUFFER
        X_ONE_INPUT_INVERTER10 N$561 OVF_SEL0 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_BUFFER3 N$577 PRE_F_0 VDD VSS ONE_INPUT_BUFFER
        X_FOUR_INPUT_AND1 N$615 N$111 N$115 N$103 N$119 N$123 N$282 VDD
+ VSS FOUR_INPUT_AND
        X_ONE_INPUT_BUFFER7 F3 N$282 VDD VSS ONE_INPUT_BUFFER
        X_ONE_INPUT_BUFFER6 F2 N$118 VDD VSS ONE_INPUT_BUFFER
        X_ONE_INPUT_BUFFER5 F1 N$103 VDD VSS ONE_INPUT_BUFFER
        X_ONE_INPUT_INVERTER3 N$629 CC1 VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_MUX1 N$475 SHIFT_OVF N$480 OVF_SEL1 N$492 VDD TWO_INPUT_MUX
        X_PROJECT_1_MUX1 N$110 N$103 N$118 N$282 A0 N$41 A1 N$31 A2 N$66
+ A3 N$20 N$40 N$30 N$65 N$19 N$577 N$36 N$70 N$26 N$577 N$36 N$70 N$26
+ N$42 N$32 N$67 N$21 N$577 N$36 N$70 N$26 N$577 N$36 N$70 N$26 A_XOR_B_0
+ N$33 N$68 A_XOR_B_2 N$287 N$288 N$289 N$159 N$287 N$288 N$289 N$159 B0
+ B1 B2 B3 N$577 N$36 N$70 N$26 CC0 N$583 CC1 N$629 CC2 N$555 CC3 N$553
+ N$287 N$288 N$289 N$159 N$287 N$288 N$289 N$159 VDD VSS VSS VSS VSS PROJECT_1_MUX
        X_ONE_INPUT_INVERTER8 N$583 CC0 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_INVERTER1 N$553 CC3 VDD VSS ONE_INPUT_INVERTER
        X_I$4 N$40 N$41 N$42 A_XOR_B_0 COUT_0 PRE_F_0 A0 ADD B0 BIN_CIN
+ CC0 N$583 CC1 N$629 CC3 N$553 VDD VSS ONE_BIT_ALU
        X_ONE_INPUT_INVERTER4 N$111 N$110 VDD VSS ONE_INPUT_INVERTER
        X_ONE_INPUT_BUFFER10 BOUT_COUT N$369 VDD VSS ONE_INPUT_BUFFER
        X_ONE_INPUT_BUFFER4 F0 N$110 VDD VSS ONE_INPUT_BUFFER
        X_ONE_INPUT_INVERTER9 N$367 N$369 VDD VSS ONE_INPUT_INVERTER
        X_TWO_INPUT_MUX2 N$480 ADD_OVF VSS OVF_SEL0 N$561 VDD TWO_INPUT_MUX
        X_SHIFTS1 N$287 N$288 N$289 N$159 SHIFT_OVF A0 A1 A2 A3 SHIFT_C_OUT
+ CC0 N$583 CC1 N$629 VDD VSS SHIFTS
        X_TWO_INPUT_AND2 ADD VDD CC0 N$583 VDD TWO_INPUT_AND
        X_ONE_INPUT_BUFFER2 COUT_2 N$568 VDD VSS ONE_INPUT_BUFFER
*
.end
