* Component: /home/ece_lab/mentor/ECE4500/HW4/function_hw4  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/HW4/function_hw4/eldonet/function_hw4_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 800N 0N 100N

* --- Waveform Outputs
.PROBE TRAN V(A) V(ANOT) V(B) V(BNOT) V(C) V(CNOT) V(F)

* --- Params
.TEMP 27

* --- Forces
VFORCE__A A VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00001111 R
VFORCE__ANOT ANOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 11110000 R
VFORCE__C C VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 01010101 R
VFORCE__CNOT CNOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 10101010 R
VFORCE__B B VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00110011 R
VFORCE__BNOT BNOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 11001100 R

* --- Libsetup

