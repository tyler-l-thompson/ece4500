* Component: /home/ece_lab/mentor/ECE4500/Project1/two_input_and/two_input_and  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/Project1/two_input_and/two_input_and/eldonet/two_input_and_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 400N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A_NOT) V(B_NOT) V(F)

* --- Params
.TEMP 27

* --- Forces
VFORCE__A_not A_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1100 R
VFORCE__B_not B_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1010 R

* --- Libsetup

