* Component: /home/ece_lab/mentor/ECE4500/HW6/npcmos_hw6  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/HW6/npcmos_hw6/eldonet/npcmos_hw6_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 1600N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A) V(B) V(C_NOT) V(CLK) V(CLK_NOT) V(F)

* --- Params
.TEMP 27

* --- Forces
VFORCE__CLK CLK VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0101010101010101 R
VFORCE__CLK_not CLK_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1010101010101010 R
VFORCE__A A VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0000000011111111 R
VFORCE__B B VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0000111100001111 R
VFORCE__C_not C_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1100110011001100 R

* --- Libsetup

