*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Tue Sep 18 2018 at 16:52:25

*
* Globals.
*
.global VSS VDD

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/HW2/HW2
*
        V2 IN VSS DC 2.5V
        V1 VDD VSS DC 2.5V
        M2 OUT IN VSS VSS NMOS L=1.2u W=2.1u M=1
        M1 OUT IN VDD VDD PMOS L=1.2u W=7.5u M=1
*
.end
