* Component: /home/ece_lab/mentor/ECE4500/Lab7/three_input_and  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/Lab7/three_input_and/eldonet/three_input_and_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 800N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A) V(B) V(C) V(F)

* --- Params
.TEMP 27

* --- Forces
VFORCE__T_3 A VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00001111 R
VFORCE__T_4 B VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00110011 R
VFORCE__T_5 C VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 01010101 R

* --- Libsetup

