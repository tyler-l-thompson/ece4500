* Component: /home/ece_lab/mentor/ECE4500/Lab7/asynchronous_sr_latch  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/Lab7/asynchronous_sr_latch/eldonet/asynchronous_sr_latch_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 800N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(CLK_18) V(CLR_NOT_18) V(QN_18) V(QN_NOT_18) V(R_18) V(S_18)

* --- Params
.TEMP 27

* --- Forces
VFORCE__CLR_not CLR_NOT_18 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00000011 R
VFORCE__R R_18 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 11100000 R
VFORCE__S S_18 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00011111 R

* --- Libsetup

