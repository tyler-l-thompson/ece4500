* Component: /home/ece_lab/mentor/4500/Project_1/Project_1_MUX  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/4500/Project_1/Project_1_MUX/eldonet/Project_1_MUX_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 1600N 0N 100N

* --- Waveform Outputs
.PROBE TRAN V(A0) V(A0_NOT) V(A1) V(A1_NOT) V(A2) V(A2_NOT) V(A3) V(A3_NOT)
+ V(A_AND_B0) V(A_AND_B1) V(A_AND_B2) V(A_AND_B3) V(A_MINUS_B0) V(A_MINUS_B1)
+ V(A_MINUS_B2) V(A_MINUS_B3) V(A_MINUS_B_WITH_BORROW0) V(A_MINUS_B_WITH_BORROW1)
+ V(A_MINUS_B_WITH_BORROW2) V(A_MINUS_B_WITH_BORROW3) V(A_OR_B0) V(A_OR_B1)
+ V(A_OR_B2) V(A_OR_B3) V(A_PLUS_B0) V(A_PLUS_B1) V(A_PLUS_B2) V(A_PLUS_B3)
+ V(A_PLUS_B_WITH_CARRY0) V(A_PLUS_B_WITH_CARRY1) V(A_PLUS_B_WITH_CARRY2)
+ V(A_PLUS_B_WITH_CARRY3) V(A_XOR_B0) V(A_XOR_B1) V(A_XOR_B2) V(A_XOR_B3) V(ASLA0)
+ V(ASLA1) V(ASLA2) V(ASLA3) V(ASRA0) V(ASRA1) V(ASRA2) V(ASRA3) V(B0) V(B1) V(B2)
+ V(B3) V(B_PLUS_ONE0) V(B_PLUS_ONE1) V(B_PLUS_ONE2) V(B_PLUS_ONE3) V(CC0)
+ V(CC0_NOT) V(CC1) V(CC1_NOT) V(CC2) V(CC2_NOT) V(CC3) V(CC3_NOT) V(F0) V(F1)
+ V(F2) V(F3) V(LSLA0) V(LSLA1) V(LSLA2) V(LSLA3) V(LSRA0) V(LSRA1) V(LSRA2)
+ V(LSRA3) V(ZERO0) V(ZERO1) V(ZERO2) V(ZERO3)

* --- Params
.TEMP 27

* --- Forces
VFORCE__A0 A0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A0_NOT A0_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1 R
VFORCE__A1 A1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A1_NOT A1_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A2 A2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A2_NOT A2_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A3_NOT A3_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A_AND_B0 A_AND_B0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A_AND_B1 A_AND_B1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1 R
VFORCE__A_AND_B2 A_AND_B2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A_AND_B3 A_AND_B3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A_MINUS_B_WITH_BORROW2 A_OR_B0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_1 A_OR_B1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_2 A_OR_B2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_3 A_OR_B3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_4 A_XOR_B0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_5 A_XOR_B1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_6 A_XOR_B2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_7 A_XOR_B3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_8 A_PLUS_B0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_9 A_PLUS_B2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_10 A_PLUS_B1 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_11 A_PLUS_B3 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_12 A_MINUS_B0 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_13 A_MINUS_B1 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_14 A_MINUS_B2 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_15 A_MINUS_B3 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_16 B0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_17 B1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_18 B2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_19 B3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_20 LSLA0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_21 LSLA1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_22 LSLA2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_23 LSLA3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_24 LSRA0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_25 LSRA1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_26 LSRA2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_27 LSRA3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_28 ASLA0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_29 ASLA1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_30 ASLA2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_31 ASLA3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_32 ASRA0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_33 ASRA1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_34 ASRA2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_35 ASRA3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_36 ZERO0 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_37 ZERO1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 0
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_38 ZERO2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_39 ZERO3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 1
+ R
VFORCE__A_MINUS_B_WITH_BORROW2_40 A_PLUS_B_WITH_CARRY0 VSS pattern 2.5 0 0 1e-12
+ 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_41 A_PLUS_B_WITH_CARRY2 VSS pattern 2.5 0 0 1e-12
+ 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_42 A_PLUS_B_WITH_CARRY3 VSS pattern 2.5 0 0 1e-12
+ 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_43 A_MINUS_B_WITH_BORROW0 VSS pattern 2.5 0 0
+ 1e-12 1e-12 1e-07 0 R
VFORCE__A_MINUS_B_WITH_BORROW2_44 A_MINUS_B_WITH_BORROW1 VSS pattern 2.5 0 0
+ 1e-12 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_45 A_MINUS_B_WITH_BORROW2 VSS pattern 2.5 0 0
+ 1e-12 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_46 A_MINUS_B_WITH_BORROW3 VSS pattern 2.5 0 0
+ 1e-12 1e-12 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_47 CC0_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 1010101010101010 R
VFORCE__A_MINUS_B_WITH_BORROW2_48 B_PLUS_ONE1 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_49 B_PLUS_ONE2 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_50 B_PLUS_ONE3 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_51 CC1 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 0011001100110011 R
VFORCE__A_MINUS_B_WITH_BORROW2_52 B_PLUS_ONE0 VSS pattern 2.5 0 0 1e-12 1e-12
+ 1e-07 1 R
VFORCE__A_MINUS_B_WITH_BORROW2_53 CC1_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 1100110011001100 R
VFORCE__A_MINUS_B_WITH_BORROW2_54 CC2 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 0000111100001111 R
VFORCE__A_MINUS_B_WITH_BORROW2_55 CC2_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 1111000011110000 R
VFORCE__A_MINUS_B_WITH_BORROW2_56 CC3 VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 0000000011111111 R
VFORCE__A_MINUS_B_WITH_BORROW2_57 CC3_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07
+ 1111111100000000 R

* --- Libsetup

