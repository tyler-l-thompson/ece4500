*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Tue Oct 30 2018 at 12:39:22

*
* Globals.
*
.global VDD VSS

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/Lab8/sense_amp/sense_amp
*
        M1 N$37 N$47 VDD VDD PMOS L=2.4u W=7.6u M=1
        V1 VDD VSS DC 2.5V
        M6 DOUTN_18 N$37 VDD VDD PMOS L=1.2u W=6.75u M=1
        M7 DOUTN_18 N$37 VSS VSS NMOS L=1.2u W=2.25u M=1
        M5 N$48 SE_18 VSS VSS NMOS L=1.2u W=2.4u M=1
        M4 N$47 DN_NOT_18 N$48 VSS NMOS L=1.2u W=2.4u M=1
        M3 N$37 DN_18 N$48 VSS NMOS L=1.2u W=2.4u M=1
        M2 N$47 N$47 VDD VDD PMOS L=2.4u W=7.6u M=1
*
.end
