* Component: /home/ece_lab/mentor/ECE4500/Project1/one_input_buffer/one_input_buffer  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/Project1/one_input_buffer/one_input_buffer/eldonet/one_input_buffer_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 200N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(IN) V(OUT)

* --- Params
.TEMP 27

* --- Forces
VFORCE__IN IN VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 01 R

* --- Libsetup

