*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Tue Oct 30 2018 at 11:35:59

*
* Globals.
*
.global VSS VDD

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/Lab8/SRAM_cell/SRAM_cell
*
        V1 VDD VSS DC 2.5V
        M5 CN_NOT_18 ROWN_18 QNOT VSS NMOS L=1.2u W=2.4u M=1
        M6 CN_18 ROWN_18 Q VSS NMOS L=1.2u W=2.4u M=1
        M1 QNOT Q VSS VSS NMOS L=1.2u W=3.0u M=1
        M2 QNOT Q VDD VDD PMOS L=1.2u W=7.8u M=1
        M3 Q QNOT VSS VSS NMOS L=1.2u W=3.0u M=1
        M4 Q QNOT VDD VDD PMOS L=1.2u W=7.8u M=1
*
.end
