* Component: /home/ece_lab/mentor/ECE4500/HW5  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/HW5/eldonet/HW5_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 800N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A) V(B) V(CNOT) V(F)

* --- Forces
VFORCE__A A VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00001111 R
VFORCE__B B VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00110011 R
VFORCE__CNOT CNOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 10101010 R

* --- Libsetup

