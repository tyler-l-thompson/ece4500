*
* .CONNECT statements
*
.CONNECT VSS 0


<<<<<<< HEAD
* ELDO netlist generated with ICnet by 'ece_lab' on Wed Sep 19 2018 at 10:47:02
=======
<<<<<<< HEAD
* ELDO netlist generated with ICnet by 'ece_lab' on Wed Sep 19 2018 at 10:47:02
=======
* ELDO netlist generated with ICnet by 'ece_lab' on Tue Sep 18 2018 at 16:52:25
>>>>>>> 559099fafff1d2d3bda55f28cce54ae15be693ac
>>>>>>> eba9bbe16f1a19bb044a525d797ef239c37b2ce1

*
* Globals.
*
.global VSS VDD

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/HW2/HW2
*
        V2 IN VSS DC 2.5V
        V1 VDD VSS DC 2.5V
        M2 OUT IN VSS VSS NMOS L=1.2u W=2.1u M=1
        M1 OUT IN VDD VDD PMOS L=1.2u W=7.5u M=1
*
.end
