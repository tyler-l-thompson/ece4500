*
* .CONNECT statements
*
.CONNECT VSS 0


* ELDO netlist generated with ICnet by 'ece_lab' on Thu Oct  4 2018 at 09:49:13

*
* Globals.
*
.global VDD VSS


*
* Component pathname : $MGC_DESIGN_KIT/symbols/ncap [SPICE]
*
*       .include /mgc/v9.0d_rhelx86linux/icstation_home/mgc_icstd_lib/mit0.25/symbols/ncap/NCAP

*
* MAIN CELL: Component pathname : /home/ece_lab/mentor/ECE4500/HW4/function_hw4
*
        X1 F VSS VSS NCAP CAPACITANCE=20F
        M10 F A N$50 VDD PMOS L=1.2u W=2.4u M=1
        M9 F ANOT N$50 VSS NMOS L=1.2u W=2.4u M=1
        M8 N$106 ANOT A VSS NMOS L=1.2u W=2.4u M=1
        M7 N$106 B A VDD PMOS L=1.2u W=2.4u M=1
        M6 N$106 BNOT A VSS NMOS L=1.2u W=2.0u M=1
        M5 BNOT B N$106 VSS NMOS L=1.2u W=2.0u M=1
        M11 F A N$106 VSS NMOS L=1.2u W=2.4u M=1
        V1 VDD VSS DC 2.5V
        M12 F ANOT N$106 VDD PMOS L=1.2u W=2.4u M=1
        M4 N$50 A ANOT VSS NMOS L=1.2u W=2.4u M=1
        M3 N$50 CNOT ANOT VDD PMOS L=1.2u W=2.4u M=1
        M2 N$50 C ANOT VSS NMOS L=1.2u W=2.0u M=1
        M1 C CNOT N$50 VSS NMOS L=1.2u W=2.0u M=1
*
.end
