* Component: /home/ece_lab/mentor/ECE4500/Project1/three_input_and/three_input_and  Viewpoint: eldonet
.INCLUDE /home/ece_lab/mentor/ECE4500/Project1/three_input_and/three_input_and/eldonet/three_input_and_eldonet.spi
.INCLUDE /home/ece_lab/mentor/mgc/mit_0.25.lib
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 800N 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A) V(B) V(B_NOT) V(C) V(C_NOT) V(F)

* --- Params
.TEMP 27

* --- Forces
VFORCE__A A VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00001111 R
VFORCE__B B VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 00110011 R
VFORCE__B_not B_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 11001100 R
VFORCE__C C VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 01010101 R
VFORCE__C_not C_NOT VSS pattern 2.5 0 0 1e-12 1e-12 1e-07 10101010 R

* --- Libsetup

